module memory(output busy, output [31:0] data_out, input clk, read_write, enable, input[1:0] access_size, input [31:0] data_in, address);

endmodule

